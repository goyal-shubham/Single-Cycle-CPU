module AndGate ( input1 , input2 , AndOut);
input input1 , input2;
output AndOut;
assign AndOut = input1 & input2;
endmodule
